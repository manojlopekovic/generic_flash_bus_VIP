/*-----------------------------------------------------------------
File name     : gfb_types defines.sv
Owner         : Manojlo Pekovic - manojlop@veriests.com
Description   : Types, enums, defines
Notes         : 
Date          : 18.03.2023.
-----------------------------------------------------------------*/
