/*-----------------------------------------------------------------
File name     : clk_types_defines.sv
Owner         : Manojlo Pekovic - manojlop@veriests.com
Description   : File that holds all enums, types and defines
Notes         : 
Date          : 12.09.2023.
-------------------------------------------------------------------
Copyright Veriest 
-----------------------------------------------------------------*/

typedef enum bit {STOP = 1'b0, START_CLK = 1'b1} t_Command;
