/*-----------------------------------------------------------------
File name     : _types_defines.sv
Owner         : Manojlo Pekovic - manojlop@veriests.com
Description   : File that holds all enums, types and defines
Notes         : 
Date          : 29.08.2023.
-------------------------------------------------------------------
Copyright Veriest 
-----------------------------------------------------------------*/
